`define GRID_SIZE 10 
`define TEST_GENERATIONS 10 
