evolve3 e0_0 (grid_evolve[0], grid[10], grid[1], grid[11], grid[0]);
evolve5 e1_0 (grid_evolve[1], grid[0], grid[10], grid[11], grid[2], grid[12], grid[1]);
evolve5 e2_0 (grid_evolve[2], grid[1], grid[11], grid[12], grid[3], grid[13], grid[2]);
evolve5 e3_0 (grid_evolve[3], grid[2], grid[12], grid[13], grid[4], grid[14], grid[3]);
evolve5 e4_0 (grid_evolve[4], grid[3], grid[13], grid[14], grid[5], grid[15], grid[4]);
evolve5 e5_0 (grid_evolve[5], grid[4], grid[14], grid[15], grid[6], grid[16], grid[5]);
evolve5 e6_0 (grid_evolve[6], grid[5], grid[15], grid[16], grid[7], grid[17], grid[6]);
evolve5 e7_0 (grid_evolve[7], grid[6], grid[16], grid[17], grid[8], grid[18], grid[7]);
evolve5 e8_0 (grid_evolve[8], grid[7], grid[17], grid[18], grid[9], grid[19], grid[8]);
evolve3 e9_0 (grid_evolve[9], grid[8], grid[18], grid[19], grid[9]);

evolve5 e0_1 (grid_evolve[10], grid[0], grid[20], grid[1], grid[11], grid[21], grid[10]);
evolve8 e1_1 (grid_evolve[11], grid[0], grid[10], grid[20], grid[1], grid[21], grid[2], grid[12], grid[22], grid[11]);
evolve8 e2_1 (grid_evolve[12], grid[1], grid[11], grid[21], grid[2], grid[22], grid[3], grid[13], grid[23], grid[12]);
evolve8 e3_1 (grid_evolve[13], grid[2], grid[12], grid[22], grid[3], grid[23], grid[4], grid[14], grid[24], grid[13]);
evolve8 e4_1 (grid_evolve[14], grid[3], grid[13], grid[23], grid[4], grid[24], grid[5], grid[15], grid[25], grid[14]);
evolve8 e5_1 (grid_evolve[15], grid[4], grid[14], grid[24], grid[5], grid[25], grid[6], grid[16], grid[26], grid[15]);
evolve8 e6_1 (grid_evolve[16], grid[5], grid[15], grid[25], grid[6], grid[26], grid[7], grid[17], grid[27], grid[16]);
evolve8 e7_1 (grid_evolve[17], grid[6], grid[16], grid[26], grid[7], grid[27], grid[8], grid[18], grid[28], grid[17]);
evolve8 e8_1 (grid_evolve[18], grid[7], grid[17], grid[27], grid[8], grid[28], grid[9], grid[19], grid[29], grid[18]);
evolve5 e9_1 (grid_evolve[19], grid[8], grid[18], grid[28], grid[9], grid[29], grid[19]);

evolve5 e0_2 (grid_evolve[20], grid[10], grid[30], grid[11], grid[21], grid[31], grid[20]);
evolve8 e1_2 (grid_evolve[21], grid[10], grid[20], grid[30], grid[11], grid[31], grid[12], grid[22], grid[32], grid[21]);
evolve8 e2_2 (grid_evolve[22], grid[11], grid[21], grid[31], grid[12], grid[32], grid[13], grid[23], grid[33], grid[22]);
evolve8 e3_2 (grid_evolve[23], grid[12], grid[22], grid[32], grid[13], grid[33], grid[14], grid[24], grid[34], grid[23]);
evolve8 e4_2 (grid_evolve[24], grid[13], grid[23], grid[33], grid[14], grid[34], grid[15], grid[25], grid[35], grid[24]);
evolve8 e5_2 (grid_evolve[25], grid[14], grid[24], grid[34], grid[15], grid[35], grid[16], grid[26], grid[36], grid[25]);
evolve8 e6_2 (grid_evolve[26], grid[15], grid[25], grid[35], grid[16], grid[36], grid[17], grid[27], grid[37], grid[26]);
evolve8 e7_2 (grid_evolve[27], grid[16], grid[26], grid[36], grid[17], grid[37], grid[18], grid[28], grid[38], grid[27]);
evolve8 e8_2 (grid_evolve[28], grid[17], grid[27], grid[37], grid[18], grid[38], grid[19], grid[29], grid[39], grid[28]);
evolve5 e9_2 (grid_evolve[29], grid[18], grid[28], grid[38], grid[19], grid[39], grid[29]);

evolve5 e0_3 (grid_evolve[30], grid[20], grid[40], grid[21], grid[31], grid[41], grid[30]);
evolve8 e1_3 (grid_evolve[31], grid[20], grid[30], grid[40], grid[21], grid[41], grid[22], grid[32], grid[42], grid[31]);
evolve8 e2_3 (grid_evolve[32], grid[21], grid[31], grid[41], grid[22], grid[42], grid[23], grid[33], grid[43], grid[32]);
evolve8 e3_3 (grid_evolve[33], grid[22], grid[32], grid[42], grid[23], grid[43], grid[24], grid[34], grid[44], grid[33]);
evolve8 e4_3 (grid_evolve[34], grid[23], grid[33], grid[43], grid[24], grid[44], grid[25], grid[35], grid[45], grid[34]);
evolve8 e5_3 (grid_evolve[35], grid[24], grid[34], grid[44], grid[25], grid[45], grid[26], grid[36], grid[46], grid[35]);
evolve8 e6_3 (grid_evolve[36], grid[25], grid[35], grid[45], grid[26], grid[46], grid[27], grid[37], grid[47], grid[36]);
evolve8 e7_3 (grid_evolve[37], grid[26], grid[36], grid[46], grid[27], grid[47], grid[28], grid[38], grid[48], grid[37]);
evolve8 e8_3 (grid_evolve[38], grid[27], grid[37], grid[47], grid[28], grid[48], grid[29], grid[39], grid[49], grid[38]);
evolve5 e9_3 (grid_evolve[39], grid[28], grid[38], grid[48], grid[29], grid[49], grid[39]);

evolve5 e0_4 (grid_evolve[40], grid[30], grid[50], grid[31], grid[41], grid[51], grid[40]);
evolve8 e1_4 (grid_evolve[41], grid[30], grid[40], grid[50], grid[31], grid[51], grid[32], grid[42], grid[52], grid[41]);
evolve8 e2_4 (grid_evolve[42], grid[31], grid[41], grid[51], grid[32], grid[52], grid[33], grid[43], grid[53], grid[42]);
evolve8 e3_4 (grid_evolve[43], grid[32], grid[42], grid[52], grid[33], grid[53], grid[34], grid[44], grid[54], grid[43]);
evolve8 e4_4 (grid_evolve[44], grid[33], grid[43], grid[53], grid[34], grid[54], grid[35], grid[45], grid[55], grid[44]);
evolve8 e5_4 (grid_evolve[45], grid[34], grid[44], grid[54], grid[35], grid[55], grid[36], grid[46], grid[56], grid[45]);
evolve8 e6_4 (grid_evolve[46], grid[35], grid[45], grid[55], grid[36], grid[56], grid[37], grid[47], grid[57], grid[46]);
evolve8 e7_4 (grid_evolve[47], grid[36], grid[46], grid[56], grid[37], grid[57], grid[38], grid[48], grid[58], grid[47]);
evolve8 e8_4 (grid_evolve[48], grid[37], grid[47], grid[57], grid[38], grid[58], grid[39], grid[49], grid[59], grid[48]);
evolve5 e9_4 (grid_evolve[49], grid[38], grid[48], grid[58], grid[39], grid[59], grid[49]);

evolve5 e0_5 (grid_evolve[50], grid[40], grid[60], grid[41], grid[51], grid[61], grid[50]);
evolve8 e1_5 (grid_evolve[51], grid[40], grid[50], grid[60], grid[41], grid[61], grid[42], grid[52], grid[62], grid[51]);
evolve8 e2_5 (grid_evolve[52], grid[41], grid[51], grid[61], grid[42], grid[62], grid[43], grid[53], grid[63], grid[52]);
evolve8 e3_5 (grid_evolve[53], grid[42], grid[52], grid[62], grid[43], grid[63], grid[44], grid[54], grid[64], grid[53]);
evolve8 e4_5 (grid_evolve[54], grid[43], grid[53], grid[63], grid[44], grid[64], grid[45], grid[55], grid[65], grid[54]);
evolve8 e5_5 (grid_evolve[55], grid[44], grid[54], grid[64], grid[45], grid[65], grid[46], grid[56], grid[66], grid[55]);
evolve8 e6_5 (grid_evolve[56], grid[45], grid[55], grid[65], grid[46], grid[66], grid[47], grid[57], grid[67], grid[56]);
evolve8 e7_5 (grid_evolve[57], grid[46], grid[56], grid[66], grid[47], grid[67], grid[48], grid[58], grid[68], grid[57]);
evolve8 e8_5 (grid_evolve[58], grid[47], grid[57], grid[67], grid[48], grid[68], grid[49], grid[59], grid[69], grid[58]);
evolve5 e9_5 (grid_evolve[59], grid[48], grid[58], grid[68], grid[49], grid[69], grid[59]);

evolve5 e0_6 (grid_evolve[60], grid[50], grid[70], grid[51], grid[61], grid[71], grid[60]);
evolve8 e1_6 (grid_evolve[61], grid[50], grid[60], grid[70], grid[51], grid[71], grid[52], grid[62], grid[72], grid[61]);
evolve8 e2_6 (grid_evolve[62], grid[51], grid[61], grid[71], grid[52], grid[72], grid[53], grid[63], grid[73], grid[62]);
evolve8 e3_6 (grid_evolve[63], grid[52], grid[62], grid[72], grid[53], grid[73], grid[54], grid[64], grid[74], grid[63]);
evolve8 e4_6 (grid_evolve[64], grid[53], grid[63], grid[73], grid[54], grid[74], grid[55], grid[65], grid[75], grid[64]);
evolve8 e5_6 (grid_evolve[65], grid[54], grid[64], grid[74], grid[55], grid[75], grid[56], grid[66], grid[76], grid[65]);
evolve8 e6_6 (grid_evolve[66], grid[55], grid[65], grid[75], grid[56], grid[76], grid[57], grid[67], grid[77], grid[66]);
evolve8 e7_6 (grid_evolve[67], grid[56], grid[66], grid[76], grid[57], grid[77], grid[58], grid[68], grid[78], grid[67]);
evolve8 e8_6 (grid_evolve[68], grid[57], grid[67], grid[77], grid[58], grid[78], grid[59], grid[69], grid[79], grid[68]);
evolve5 e9_6 (grid_evolve[69], grid[58], grid[68], grid[78], grid[59], grid[79], grid[69]);

evolve5 e0_7 (grid_evolve[70], grid[60], grid[80], grid[61], grid[71], grid[81], grid[70]);
evolve8 e1_7 (grid_evolve[71], grid[60], grid[70], grid[80], grid[61], grid[81], grid[62], grid[72], grid[82], grid[71]);
evolve8 e2_7 (grid_evolve[72], grid[61], grid[71], grid[81], grid[62], grid[82], grid[63], grid[73], grid[83], grid[72]);
evolve8 e3_7 (grid_evolve[73], grid[62], grid[72], grid[82], grid[63], grid[83], grid[64], grid[74], grid[84], grid[73]);
evolve8 e4_7 (grid_evolve[74], grid[63], grid[73], grid[83], grid[64], grid[84], grid[65], grid[75], grid[85], grid[74]);
evolve8 e5_7 (grid_evolve[75], grid[64], grid[74], grid[84], grid[65], grid[85], grid[66], grid[76], grid[86], grid[75]);
evolve8 e6_7 (grid_evolve[76], grid[65], grid[75], grid[85], grid[66], grid[86], grid[67], grid[77], grid[87], grid[76]);
evolve8 e7_7 (grid_evolve[77], grid[66], grid[76], grid[86], grid[67], grid[87], grid[68], grid[78], grid[88], grid[77]);
evolve8 e8_7 (grid_evolve[78], grid[67], grid[77], grid[87], grid[68], grid[88], grid[69], grid[79], grid[89], grid[78]);
evolve5 e9_7 (grid_evolve[79], grid[68], grid[78], grid[88], grid[69], grid[89], grid[79]);

evolve5 e0_8 (grid_evolve[80], grid[70], grid[90], grid[71], grid[81], grid[91], grid[80]);
evolve8 e1_8 (grid_evolve[81], grid[70], grid[80], grid[90], grid[71], grid[91], grid[72], grid[82], grid[92], grid[81]);
evolve8 e2_8 (grid_evolve[82], grid[71], grid[81], grid[91], grid[72], grid[92], grid[73], grid[83], grid[93], grid[82]);
evolve8 e3_8 (grid_evolve[83], grid[72], grid[82], grid[92], grid[73], grid[93], grid[74], grid[84], grid[94], grid[83]);
evolve8 e4_8 (grid_evolve[84], grid[73], grid[83], grid[93], grid[74], grid[94], grid[75], grid[85], grid[95], grid[84]);
evolve8 e5_8 (grid_evolve[85], grid[74], grid[84], grid[94], grid[75], grid[95], grid[76], grid[86], grid[96], grid[85]);
evolve8 e6_8 (grid_evolve[86], grid[75], grid[85], grid[95], grid[76], grid[96], grid[77], grid[87], grid[97], grid[86]);
evolve8 e7_8 (grid_evolve[87], grid[76], grid[86], grid[96], grid[77], grid[97], grid[78], grid[88], grid[98], grid[87]);
evolve8 e8_8 (grid_evolve[88], grid[77], grid[87], grid[97], grid[78], grid[98], grid[79], grid[89], grid[99], grid[88]);
evolve5 e9_8 (grid_evolve[89], grid[78], grid[88], grid[98], grid[79], grid[99], grid[89]);

evolve3 e0_9 (grid_evolve[90], grid[80], grid[81], grid[91], grid[90]);
evolve5 e1_9 (grid_evolve[91], grid[80], grid[90], grid[81], grid[82], grid[92], grid[91]);
evolve5 e2_9 (grid_evolve[92], grid[81], grid[91], grid[82], grid[83], grid[93], grid[92]);
evolve5 e3_9 (grid_evolve[93], grid[82], grid[92], grid[83], grid[84], grid[94], grid[93]);
evolve5 e4_9 (grid_evolve[94], grid[83], grid[93], grid[84], grid[85], grid[95], grid[94]);
evolve5 e5_9 (grid_evolve[95], grid[84], grid[94], grid[85], grid[86], grid[96], grid[95]);
evolve5 e6_9 (grid_evolve[96], grid[85], grid[95], grid[86], grid[87], grid[97], grid[96]);
evolve5 e7_9 (grid_evolve[97], grid[86], grid[96], grid[87], grid[88], grid[98], grid[97]);
evolve5 e8_9 (grid_evolve[98], grid[87], grid[97], grid[88], grid[89], grid[99], grid[98]);
evolve3 e9_9 (grid_evolve[99], grid[88], grid[98], grid[89], grid[99]);

